
module music_ROM(
	input clk,
	input [7:0] address,
	output reg [7:0] note
);

always @(posedge clk)
case(address)

//Oh dont you dare...
      0: note<= 8'd31;  //D
      1: note<= 8'd31;  //D
	  2: note<= 8'd31;  //D
	  3: note<= 8'd31;  //D
	  4: note<= 8'd31;  //D
	  5: note<= 8'd31;  //D
      
      6: note<= 8'd31;  //D
      7: note<= 8'd31;  //D
      8: note<= 8'd31;  //D
      9: note<= 8'd31;  //D
      10: note<= 8'd31;  //D
      11: note<= 8'd31;  //D
      
      //Just keep your eyes....
      12: note<= 8'd31;  //D
	  13: note<= 8'd31;  //D
	  14: note<= 8'd31;  //D
	  15: note<= 8'd31;  //D
	  16: note<= 8'd31;  //D      
	  17: note<= 8'd31;  //D 
      
      18: note<= 8'd31;  //D 
      19: note<= 8'd31;  //D 
      20: note<= 8'd31;  //D 
      21: note<= 8'd31;  //D 
      22: note<= 8'd21;  //Eb
      23: note<= 8'd21;  //Eb

      //I said youre holding back....
      24: note<= 8'd31;  //D
	  25: note<= 8'd31;  //D
	  26: note<= 8'd31;  //D
	  27: note<= 8'd31;  //D
	  28: note<= 8'd31;  //D
	  29: note<= 8'd31;  //D
      
      30: note<= 8'd31;  //D
      31: note<= 8'd31;  //D
      32: note<= 8'd31;  //D
      33: note<= 8'd31;  //D
      34: note<= 8'd31;  //D
      35: note<= 8'd31;  //D
      
      //She said shut up.,...
      36: note<= 8'd31;  //D
	  37: note<= 8'd31;  //D
      38: note<= 8'd31;  //D
	  39: note<= 8'd31;  //D
      
      40: note<= 8'd25;  //Ab
      41: note<= 8'd25;  //Ab
      
      42: note<= 8'd25;  //Ab
      43: note<= 8'd25;  //Ab
      
      44: note<= 8'd23;  //F
      45: note<= 8'd23;  //F
      
      46: note<= 8'd21; //Eb
      47: note<= 8'd21; //Eb
      
      48: note<= 8'd31;  //D
      49: note<= 8'd31;  //D
      
      50:  note<= 8'd31;  //D
      51: note<= 8'd31;  //D
      
      //This woman is my ....
      52: note<= 8'd31;  //D
      53: note<= 8'd31;  //D
      
      54: note<= 8'd28; //Bb
      55: note<= 8'd28; //Bb
      
      56: note<= 8'd31; //D
      57: note<= 8'd31; //D
      
      58: note<= 8'd31; //D
      59: note<= 8'd31; //D
      
      60: note<= 8'd21; //Eb
      61: note<= 8'd21; //Eb
      
      62: note<= 8'd23; //F
      63: note<= 8'd23; //F
      
      64: note<= 8'd31; //D
      65: note<= 8'd31; //D
      
      66: note<= 8'd21; //Eb
      67: note<= 8'd21; //Eb

//She siad ohh oh
      68: note<= 8'd31; //D
      69: note<= 8'd31; //D
      
      70: note<= 8'd31; //D
      71: note<= 8'd31; //D
      
      72: note<= 8'd25; //Ab
      73: note<= 8'd25; //Ab
      
      74: note<= 8'd23; //F
      75: note<= 8'd23; //F
      
      76: note<= 8'd28;  //Bb
      77: note<= 8'd28;  //Bb
      
      //Shut up and dance...
      78: note<= 8'd26; //Ab
      79: note<= 8'd26; //Ab
      
      80: note<= 8'd26; //Ab
      81: note<= 8'd26; //Ab
      
      82: note<= 8'd23; //F
      83: note<= 8'd23; //F
      
      84: note<= 8'd21; //Eb
      85: note<= 8'd21; //Eb
      
      86: note<= 8'd31;  //D
      87: note <= 8'd31;    //D
      
      88: note<= 8'd31;  //D
      89: note <= 8'd31;    //D
      
      //We were victims of the night
      90: note<= 8'd31; //D
      91: note<= 8'd31; //D
      
      92: note<= 8'd31; //D
	  93: note<= 8'd31; //D
      
      94: note<= 8'd31;  //D
      95: note<= 8'd31; //D
      
      96: note<= 8'd28;  //Bb
      97: note<= 8'd28;  //Bb
      
	  98: note<= 8'd26; //Ab
      100: note<= 8'd26; //Ab

      101: note<= 8'd31; //D
      102: note<= 8'd31; //D
      
      //FIX THIS SHIT :)))))))
      
      /*
//The chemical, physical,.....
	  50: note<= 8'd31;  //D
	  51: note<= 8'd31;  //D
	  52: note<= 8'd31;  //D
	  53: note<= 8'd28;  //Bb
	  54: note<= 8'd31;  //D
	  55: note<= 8'd31;  //D
	  56: note<= 8'd28;  //Bb	 
      57: note<= 8'd31;  //D
      58: note<= 8'd21;  //Eb
      59: note<= 8'd23;   //F

      //Helpless to the bass....
      60: note<= 8'd31;   //D
	  61: note<= 8'd31;   //D
	  62: note<= 8'd31;   //D   
	  63: note<= 8'd28;   //Bb
	  64: note<= 8'd31;   //D
	  65: note<= 8'd28;   //Bb
	  66: note<= 8'd26;   //Ab
	  67: note<= 8'd28;   //Bb
	  68: note<= 8'd31;   //D
	 
     //Oh we were bound
     69: note<= 8'd31;   //D
	  70: note<= 8'd31;   //D
	  71: note<= 8'd31;   //D
	  72: note<= 8'd26;   //Ab
	  73: note<= 8'd23;   //F
	  74: note<= 8'd23;   //F
	  75: note<= 8'd21;   //Eb
	  76: note<= 8'd21;   //Eb
	  77: note<= 8'd31;   //D
	 
     //Bound to get
      78: note<= 8'd26;    //Ab
	  79: note<= 8'd23;    //F
	  80: note<= 8'd23;    //F
	  81: note<= 8'd21;    //Eb
	  82: note<= 8'd21;    //Eb
	  83: note<= 8'd31;    //D
      
      //She took my arm
	  84: note<= 8'd31;    //D
	  85: note<= 8'd31;    //D
	  86: note<= 8'd21;    //Eb
	  87: note<= 8'd21;    //Eb
      
      //I dont know how it...
	  88: note<= 8'd23;   //F
	  89: note<= 8'd23;   //F
	 90: note<= 8'd23;   //F 
	 91: note<= 8'd24;   //Gb
	 92: note<= 8'd23;   //F
	 93: note<= 8'd21;   //Eb
	 94: note<= 8'd31;   //D
	
    //We took the floor...
     95: note<= 8'd31;  //D
	 96: note<= 8'd31;  //D
	 97: note<= 8'd21;  //Eb
	 98: note<= 8'd21;  //Eb
	 99: note<= 8'd31;  //D
	 100: note<= 8'd31;  //D
	 101: note<= 8'd26;  //Ab
	
    //Oh dont you dare
     102: note<= 8'd31;  //D
	 103: note<= 8'd31;  //D
	 104: note<= 8'd31;  //D
	 105: note<= 8'd31;  //D
	 106: note<= 8'd31;  //D
	 107: note<= 8'd31;  //D
     
     //Just keep
	 108: note<= 8'd31;  //D
	 109: note<= 8'd31;  //D
	 110: note<= 8'd31;  //D
	 111: note<= 8'd31;  //D
	 112: note<= 8'd31;  //D
	 113: note<= 8'd21; //Eb
     
     //I said youre holding
	 114: note<= 8'd31;  //D
	 115: note<= 8'd31;  //D
	 116: note<= 8'd31;  //D
	 117: note<= 8'd31;  //D
	 118: note<= 8'd31;  //D
	 119: note<= 8'd31;  //D
     
     //She said Shut up and dance
	 120: note<= 8'd31;  //D
	 121: note<= 8'd31;  //D
	 122: note<= 8'd26;  //Ab
	 123: note<= 8'd26;  //Ab
	 124: note<= 8'd23;   //F 
	 125: note<= 8'd21; //Eb
	 126: note<= 8'd31;  //D
	 127: note<= 8'd31;  //D
     
     //This woman is my destiny
      128: note<= 8'd31;  //D
      129: note<= 8'd28; //Bb
      130: note<= 8'd31; //D
      131: note<= 8'd31; //D
      132: note<= 8'd21; //Eb
      133: note<= 8'd23; //F
      134: note<= 8'd31; //D
      135: note<= 8'd21; //Eb
     
      //She said Oh oh oh
      136: note<= 8'd31; //D
      137: note<= 8'd31; //D
      138: note<= 8'd25; //Ab
      139: note<= 8'd23; //F
      140: note<= 8'd28;  //Bb
     
     //Shut up and dance
     141: note<= 8'd31;  //D
	 142: note<= 8'd31;  //D
	 143: note<= 8'd26;  //Ab
	 144: note<= 8'd26;  //Ab
	 145: note<= 8'd23;   //F 
	 146: note<= 8'd21; //Eb
	 147: note<= 8'd31;  //D
	 148: note<= 8'd31;  //D
     
     //A backless dress
	149: note<= 8'd31;  //D
	150: note<= 8'd31;  //D
	151: note<= 8'd31;  //D
	152: note<= 8'd31;  //D
    
    //and some beat up sneaks 
	153: note<= 8'd28;  //Bb
	154: note<= 8'd26;  //Ab
	155: note<= 8'd26;  //Ab
	156: note<= 8'd28;  //Bb
	157: note<= 8'd31;  //D
   
    //My disco tech
	158: note<= 8'd31;  //D
	159: note<= 8'd31;  //D
	160: note<= 8'd31;  //D
	161: note<= 8'd28;  //Bb
	162: note<= 8'd31;  //D
	163: note<= 8'd31;  //D
	164: note<= 8'd28;  //Bb
	165: note<= 8'd31;  //D
	166: note<= 8'd21;  //Eb
	167: note<= 8'd23;  //F
    
   //I felt it.. 
	168: note<= 8'd31;  //D
	169: note<= 8'd31;  //D
	170: note<= 8'd31;  //D
	171: note<= 8'd31;  //D
	172: note<= 8'd31;  //D
	173: note<= 8'd31;  //D
	174: note<= 8'd28;  //Bb
	175: note<= 8'd26;  //Ab
	176: note<= 8'd26;  //Ab
	177: note<= 8'd28;  //Bb
	178: note<= 8'd31;  //D
    
    //I knew we...
	179: note<= 8'd31;  //D
	180: note<= 8'd31;  //D
	181: note<= 8'd31;  //D
	182: note<= 8'd31;  //D
	183: note<= 8'd26;  //Ab
	184: note<= 8'd23;  //F
	185: note<= 8'd23;  //F
	186: note<= 8'd21;  //Eb
	187: note<= 8'd21;  //Eb
	188: note<= 8'd31;  //D
    
    //Bound to be...
	189: note<= 8'd26;  //Ab
	190: note<= 8'd23;  //F
	191: note<= 8'd23;  //F
	192: note<= 8'd21;  //Eb
	193: note<= 8'd21;  //Eb
	194: note<= 8'd31;  //D

    //She took my arm
	195: note<= 8'd31;  //D
	196: note<= 8'd31;  //D
	197: note<= 8'd31;  //D
	198: note<= 8'd31;  //D
    
    //I don't know...
	199: note<= 8'd23;  //F
	200: note<= 8'd23;  //F
	201: note<= 8'd23;  //F
	202: note<= 8'd24;  //Gb
	203: note<= 8'd23;  //F
	204: note<= 8'd21;  //Eb
	205: note<= 8'd31;  //D
    
    //We took the floor...
	206: note<= 8'd31;  //D
	207: note<= 8'd31;  //D
	208: note<= 8'd21;  //Eb
	209: note<= 8'd21;  //Eb
	210: note<= 8'd31;  //D
	211: note<= 8'd31;  //D
	212: note<= 8'd31;  //D
	213: note<= 8'd26;  //Ab
    
    //Oh don't you 
	214: note<= 8'd31;  //D
	215: note<= 8'd31;  //D
	216: note<= 8'd31;  //D
	217: note<= 8'd31;  //D
	218: note<= 8'd31;  //D
	219: note<= 8'd31;  //D
    
    //I said you're...
	220: note<= 8'd31;  //D
	221: note<= 8'd31;  //D
	222: note<= 8'd31;  //D
	223: note<= 8'd31;  //D
	224: note<= 8'd31;  //D
	225: note<= 8'd31;  //D
    
    //She said, Shut up
	226: note<= 8'd31;  //D
	227: note<= 8'd31;  //D
	228: note<= 8'd26;  //Ab
	229: note<= 8'd26;  //Ab
	230: note<= 8'd23;  //F
	231: note<= 8'd21;  //Eb
	232: note<= 8'd31;   //D
	233: note<= 8'd31;  //D
    
    //This woman is....
	234: note<= 8'd31;  //D
	235: note<= 8'd28;  //Bb
	236: note<= 8'd31;  //D
	237: note<= 8'd31;  //D
	238: note<= 8'd21;  //Eb
	239: note<= 8'd23;  //F
	240: note<= 8'd31;  //D
	241: note<= 8'd21;  //Eb
    
    //She said, Oh
	242: note<= 8'd31;  //D
	243: note<= 8'd31;  //D
	244: note<= 8'd26;  //Ab
	245: note<= 8'd23;  //F
	246: note<= 8'd28;  //Bb
    
    //Shut up and...
	247: note<= 8'd26;  //Ab
	248: note<= 8'd26;  //Ab
	249: note<= 8'd23;  //F
	250: note<= 8'd21;  //Eb
	251: note<= 8'd31;  //D
	252: note<= 8'd31;  //D
      
      //Deep in her eyes
    253: note<= 8'd31;  //D
    254: note<= 8'd31;  //D
    255: note<= 8'd21;  //Eb
    256: note<= 8'd21;  //Eb
    
    //I think I see...
    257: note<= 8'd23;  //F
    258: note<= 8'd23;  //F
    259: note<= 8'd23;  //F
    260: note<= 8'd25;  //Gb
    261: note<= 8'd23;  //F
    262: note<= 8'd21;  //Eb
    263: note<= 8'd31;  //Db

    //I realize this is my ....
    264: note<= 8'd31;  //Db
    265: note<= 8'd31;  //Db
    266: note<= 8'd21;  //Eb
    267: note<= 8'd21;  //Eb
    268: note<= 8'd23;  //F
    269: note<= 8'd23;  //F
    270: note<= 8'd23;  //F
    271: note<= 8'd26;  //Ab
    272: note<= 8'd26;  //Ab

    //She took my arm
    273: note<= 8'd31;  //Db
    274: note<= 8'd31;  //Db
    275: note<= 8'd31;  //Db
    276: note<= 8'd31;  //Db

    //I dont know how it happened
	  279: note<= 8'd23;   //F
	  280: note<= 8'd23;   //F
	 281: note<= 8'd23;   //F 
	 282: note<= 8'd24;   //Gb
	 283: note<= 8'd23;   //F
	 284: note<= 8'd21;   //Eb
	 285: note<= 8'd31;   //D
     
     //We took the floor
    286: note<= 8'd31;  //D
	287: note<= 8'd31;  //D
	288: note<= 8'd21;  //Eb
	289: note<= 8'd21;  //Eb
	290: note<= 8'd31;  //D
	291: note<= 8'd31;  //D
	292: note<= 8'd31;  //D
	293: note<= 8'd26;  //Ab
     
     //Oh dont you dare
     294: note<= 8'd31;  //D
     295: note<= 8'd31;  //D
	 296: note<= 8'd31;  //D
	  297: note<= 8'd31;  //D
	  298: note<= 8'd31;  //D
	 299: note<= 8'd31;  //D
     
     //Just keep
      300: note<= 8'd31;  //D
	  301: note<= 8'd31;  //D
	  302: note<= 8'd31;  //D
	  303: note<= 8'd31;  //D
	  304: note<= 8'd31;  //D      
	  305: note<= 8'd21;  //Eb
     
 //I said youre holding back....
      306: note<= 8'd31;  //D
	  307: note<= 8'd31;  //D
	  308: note<= 8'd31;  //D
	  309: note<= 8'd31;  //D
	  310: note<= 8'd31;  //D
	  311: note<= 8'd31;  //D
      
      //She said shut up.,...
      312: note<= 8'd31;  //D
	  313: note<= 8'd31;  //D
	  314: note<= 8'd25;  //Ab
      315: note<= 8'd25;  //Ab
      316: note<= 8'd23;  //F
      317: note<= 8'd21; //Eb
      318: note<= 8'd31;  //D
      319: note<= 8'd31;  //D
      
      //This woman is my ....
      320: note<= 8'd31;  //D
      321: note<= 8'd28; //Bb
      322: note<= 8'd31; //D
      323: note<= 8'd31; //D
      324: note<= 8'd21; //Eb
      325: note<= 8'd23; //F
      326: note<= 8'd31; //D
      327: note<= 8'd21; //Eb

//She siad ohh oh
      328: note<= 8'd31; //D
      329: note<= 8'd31; //D
      330: note<= 8'd25; //Ab
      331: note<= 8'd23; //F
      332: note<= 8'd28;  //Bb
      
      //Shut up and dance...
      333: note<= 8'd26; //Ab
      334: note<= 8'd26; //Ab
      335: note<= 8'd23; //F
      336: note<= 8'd21; //Eb
      337: note<= 8'd31;  //D
      338: note <= 8'd31;    //D
*/

/*
//Oh dont you dare...
      0: note<= 8'd31;  //D
      1: note<= 8'd31;  //D
	  2: note<= 8'd31;  //D
	  3: note<= 8'd31;  //D
	  4: note<= 8'd31;  //D
	  5: note<= 8'd31;  //D
      
      //Just keep your eyes....
      6: note<= 8'd31;  //D
	  7: note<= 8'd31;  //D
	  8: note<= 8'd31;  //D
	  9: note<= 8'd31;  //D
	  10: note<= 8'd31;  //D      
	  11: note<= 8'd21;  //Eb
      
      //I said youre holding back....
      12: note<= 8'd31;  //D
	  13: note<= 8'd31;  //D
	  14: note<= 8'd31;  //D
	  15: note<= 8'd31;  //D
	  16: note<= 8'd31;  //D
	  17: note<= 8'd31;  //D
      
      //She said shut up.,...
      18: note<= 8'd31;  //D
	  19: note<= 8'd31;  //D
	  20: note<= 8'd25;  //Ab
      21: note<= 8'd25;  //Ab
      22: note<= 8'd23;  //F
      23: note<= 8'd21; //Eb
      24: note<= 8'd31;  //D
      25: note<= 8'd31;  //D
      
      //This woman is my ....
      26: note<= 8'd31;  //D
      27: note<= 8'd28; //Bb
      28: note<= 8'd31; //D
      29: note<= 8'd31; //D
      30: note<= 8'd21; //Eb
      31: note<= 8'd23; //F
      32: note<= 8'd31; //D
      33: note<= 8'd21; //Eb

//She siad ohh oh
      34: note<= 8'd31; //D
      35: note<= 8'd31; //D
      36: note<= 8'd25; //Ab
      37: note<= 8'd23; //F
      38: note<= 8'd28;  //Bb
      
      //Shut up and dance...
      39: note<= 8'd26; //Ab
      40: note<= 8'd26; //Ab
      41: note<= 8'd23; //F
      42: note<= 8'd21; //Eb
      42: note<= 8'd31;  //D
      43: note <= 8'd31;    //D
      
      //We were victims of the night
      44: note<= 8'd31; //D
      45: note<= 8'd31; //D
	  46: note<= 8'd31;  //D
      47: note<= 8'd28;  //Bb
	  48: note<= 8'd26; //Ab
      49: note<= 8'd31; //D

//The chemical, physical,.....
	  50: note<= 8'd31;  //D
	  51: note<= 8'd31;  //D
	  52: note<= 8'd31;  //D
	  53: note<= 8'd28;  //Bb
	  54: note<= 8'd31;  //D
	  55: note<= 8'd31;  //D
	  56: note<= 8'd28;  //Bb	 
      57: note<= 8'd31;  //D
      58: note<= 8'd21;  //Eb
      59: note<= 8'd23;   //F

      //Helpless to the bass....
      60: note<= 8'd31;   //D
	  61: note<= 8'd31;   //D
	  62: note<= 8'd31;   //D   
	  63: note<= 8'd28;   //Bb
	  64: note<= 8'd31;   //D
	  65: note<= 8'd28;   //Bb
	  66: note<= 8'd26;   //Ab
	  67: note<= 8'd28;   //Bb
	  68: note<= 8'd31;   //D
	 
     //Oh we were bound
     69: note<= 8'd31;   //D
	  70: note<= 8'd31;   //D
	  71: note<= 8'd31;   //D
	  72: note<= 8'd26;   //Ab
	  73: note<= 8'd23;   //F
	  74: note<= 8'd23;   //F
	  75: note<= 8'd21;   //Eb
	  76: note<= 8'd21;   //Eb
	  77: note<= 8'd31;   //D
	 
     //Bound to get
      78: note<= 8'd26;    //Ab
	  79: note<= 8'd23;    //F
	  80: note<= 8'd23;    //F
	  81: note<= 8'd21;    //Eb
	  82: note<= 8'd21;    //Eb
	  83: note<= 8'd31;    //D
      
      //She took my arm
	  84: note<= 8'd31;    //D
	  85: note<= 8'd31;    //D
	  86: note<= 8'd21;    //Eb
	  87: note<= 8'd21;    //Eb
      
      //I dont know how it...
	  88: note<= 8'd23;   //F
	  89: note<= 8'd23;   //F
	 90: note<= 8'd23;   //F 
	 91: note<= 8'd24;   //Gb
	 92: note<= 8'd23;   //F
	 93: note<= 8'd21;   //Eb
	 94: note<= 8'd31;   //D
	
    //We took the floor...
     95: note<= 8'd31;  //D
	 96: note<= 8'd31;  //D
	 97: note<= 8'd21;  //Eb
	 98: note<= 8'd21;  //Eb
	 99: note<= 8'd31;  //D
	 100: note<= 8'd31;  //D
	 101: note<= 8'd26;  //Ab
	
    //Oh dont you dare
     102: note<= 8'd31;  //D
	 103: note<= 8'd31;  //D
	 104: note<= 8'd31;  //D
	 105: note<= 8'd31;  //D
	 106: note<= 8'd31;  //D
	 107: note<= 8'd31;  //D
     
     //Just keep
	 108: note<= 8'd31;  //D
	 109: note<= 8'd31;  //D
	 110: note<= 8'd31;  //D
	 111: note<= 8'd31;  //D
	 112: note<= 8'd31;  //D
	 113: note<= 8'd21; //Eb
     
     //I said youre holding
	 114: note<= 8'd31;  //D
	 115: note<= 8'd31;  //D
	 116: note<= 8'd31;  //D
	 117: note<= 8'd31;  //D
	 118: note<= 8'd31;  //D
	 119: note<= 8'd31;  //D
     
     //She said Shut up and dance
	 120: note<= 8'd31;  //D
	 121: note<= 8'd31;  //D
	 122: note<= 8'd26;  //Ab
	 123: note<= 8'd26;  //Ab
	 124: note<= 8'd23;   //F 
	 125: note<= 8'd21; //Eb
	 126: note<= 8'd31;  //D
	 127: note<= 8'd31;  //D
     
     //This woman is my destiny
      128: note<= 8'd31;  //D
      129: note<= 8'd28; //Bb
      130: note<= 8'd31; //D
      131: note<= 8'd31; //D
      132: note<= 8'd21; //Eb
      133: note<= 8'd23; //F
      134: note<= 8'd31; //D
      135: note<= 8'd21; //Eb
     
      //She said Oh oh oh
      136: note<= 8'd31; //D
      137: note<= 8'd31; //D
      138: note<= 8'd25; //Ab
      139: note<= 8'd23; //F
      140: note<= 8'd28;  //Bb
     
     //Shut up and dance
     141: note<= 8'd31;  //D
	 142: note<= 8'd31;  //D
	 143: note<= 8'd26;  //Ab
	 144: note<= 8'd26;  //Ab
	 145: note<= 8'd23;   //F 
	 146: note<= 8'd21; //Eb
	 147: note<= 8'd31;  //D
	 148: note<= 8'd31;  //D
     
     //A backless dress
	149: note<= 8'd31;  //D
	150: note<= 8'd31;  //D
	151: note<= 8'd31;  //D
	152: note<= 8'd31;  //D
    
    //and some beat up sneaks 
	153: note<= 8'd28;  //Bb
	154: note<= 8'd26;  //Ab
	155: note<= 8'd26;  //Ab
	156: note<= 8'd28;  //Bb
	157: note<= 8'd31;  //D
   
    //My disco tech
	158: note<= 8'd31;  //D
	159: note<= 8'd31;  //D
	160: note<= 8'd31;  //D
	161: note<= 8'd28;  //Bb
	162: note<= 8'd31;  //D
	163: note<= 8'd31;  //D
	164: note<= 8'd28;  //Bb
	165: note<= 8'd31;  //D
	166: note<= 8'd21;  //Eb
	167: note<= 8'd23;  //F
    
   //I felt it.. 
	168: note<= 8'd31;  //D
	169: note<= 8'd31;  //D
	170: note<= 8'd31;  //D
	171: note<= 8'd31;  //D
	172: note<= 8'd31;  //D
	173: note<= 8'd31;  //D
	174: note<= 8'd28;  //Bb
	175: note<= 8'd26;  //Ab
	176: note<= 8'd26;  //Ab
	177: note<= 8'd28;  //Bb
	178: note<= 8'd31;  //D
    
    //I knew we...
	179: note<= 8'd31;  //D
	180: note<= 8'd31;  //D
	181: note<= 8'd31;  //D
	182: note<= 8'd31;  //D
	183: note<= 8'd26;  //Ab
	184: note<= 8'd23;  //F
	185: note<= 8'd23;  //F
	186: note<= 8'd21;  //Eb
	187: note<= 8'd21;  //Eb
	188: note<= 8'd31;  //D
    
    //Bound to be...
	189: note<= 8'd26;  //Ab
	190: note<= 8'd23;  //F
	191: note<= 8'd23;  //F
	192: note<= 8'd21;  //Eb
	193: note<= 8'd21;  //Eb
	194: note<= 8'd31;  //D

    //She took my arm
	195: note<= 8'd31;  //D
	196: note<= 8'd31;  //D
	197: note<= 8'd31;  //D
	198: note<= 8'd31;  //D
    
    //I don't know...
	199: note<= 8'd23;  //F
	200: note<= 8'd23;  //F
	201: note<= 8'd23;  //F
	202: note<= 8'd24;  //Gb
	203: note<= 8'd23;  //F
	204: note<= 8'd21;  //Eb
	205: note<= 8'd31;  //D
    
    //We took the floor...
	206: note<= 8'd31;  //D
	207: note<= 8'd31;  //D
	208: note<= 8'd21;  //Eb
	209: note<= 8'd21;  //Eb
	210: note<= 8'd31;  //D
	211: note<= 8'd31;  //D
	212: note<= 8'd31;  //D
	213: note<= 8'd26;  //Ab
    
    //Oh don't you 
	214: note<= 8'd31;  //D
	215: note<= 8'd31;  //D
	216: note<= 8'd31;  //D
	217: note<= 8'd31;  //D
	218: note<= 8'd31;  //D
	219: note<= 8'd31;  //D
    
    //I said you're...
	220: note<= 8'd31;  //D
	221: note<= 8'd31;  //D
	222: note<= 8'd31;  //D
	223: note<= 8'd31;  //D
	224: note<= 8'd31;  //D
	225: note<= 8'd31;  //D
    
    //She said, Shut up
	226: note<= 8'd31;  //D
	227: note<= 8'd31;  //D
	228: note<= 8'd26;  //Ab
	229: note<= 8'd26;  //Ab
	230: note<= 8'd23;  //F
	231: note<= 8'd21;  //Eb
	232: note<= 8'd31;   //D
	233: note<= 8'd31;  //D
    
    //This woman is....
	234: note<= 8'd31;  //D
	235: note<= 8'd28;  //Bb
	236: note<= 8'd31;  //D
	237: note<= 8'd31;  //D
	238: note<= 8'd21;  //Eb
	239: note<= 8'd23;  //F
	240: note<= 8'd31;  //D
	241: note<= 8'd21;  //Eb
    
    //She said, Oh
	242: note<= 8'd31;  //D
	243: note<= 8'd31;  //D
	244: note<= 8'd26;  //Ab
	245: note<= 8'd23;  //F
	246: note<= 8'd28;  //Bb
    
    //Shut up and...
	247: note<= 8'd26;  //Ab
	248: note<= 8'd26;  //Ab
	249: note<= 8'd23;  //F
	250: note<= 8'd21;  //Eb
	251: note<= 8'd31;  //D
	252: note<= 8'd31;  //D
      
      //Deep in her eyes
    253: note<= 8'd31;  //D
    254: note<= 8'd31;  //D
    255: note<= 8'd21;  //Eb
    256: note<= 8'd21;  //Eb
    
    //I think I see...
    257: note<= 8'd23;  //F
    258: note<= 8'd23;  //F
    259: note<= 8'd23;  //F
    260: note<= 8'd25;  //Gb
    261: note<= 8'd23;  //F
    262: note<= 8'd21;  //Eb
    263: note<= 8'd31;  //Db

    //I realize this is my ....
    264: note<= 8'd31;  //Db
    265: note<= 8'd31;  //Db
    266: note<= 8'd21;  //Eb
    267: note<= 8'd21;  //Eb
    268: note<= 8'd23;  //F
    269: note<= 8'd23;  //F
    270: note<= 8'd23;  //F
    271: note<= 8'd26;  //Ab
    272: note<= 8'd26;  //Ab

    //She took my arm
    273: note<= 8'd31;  //Db
    274: note<= 8'd31;  //Db
    275: note<= 8'd31;  //Db
    276: note<= 8'd31;  //Db

    //I dont know how it happened
	  279: note<= 8'd23;   //F
	  280: note<= 8'd23;   //F
	 281: note<= 8'd23;   //F 
	 282: note<= 8'd24;   //Gb
	 283: note<= 8'd23;   //F
	 284: note<= 8'd21;   //Eb
	 285: note<= 8'd31;   //D
     
     //We took the floor
    286: note<= 8'd31;  //D
	287: note<= 8'd31;  //D
	288: note<= 8'd21;  //Eb
	289: note<= 8'd21;  //Eb
	290: note<= 8'd31;  //D
	291: note<= 8'd31;  //D
	292: note<= 8'd31;  //D
	293: note<= 8'd26;  //Ab
     
     //Oh dont you dare
     294: note<= 8'd31;  //D
     295: note<= 8'd31;  //D
	 296: note<= 8'd31;  //D
	  297: note<= 8'd31;  //D
	  298: note<= 8'd31;  //D
	 299: note<= 8'd31;  //D
     
     //Just keep
      300: note<= 8'd31;  //D
	  301: note<= 8'd31;  //D
	  302: note<= 8'd31;  //D
	  303: note<= 8'd31;  //D
	  304: note<= 8'd31;  //D      
	  305: note<= 8'd21;  //Eb
     
 //I said youre holding back....
      306: note<= 8'd31;  //D
	  307: note<= 8'd31;  //D
	  308: note<= 8'd31;  //D
	  309: note<= 8'd31;  //D
	  310: note<= 8'd31;  //D
	  311: note<= 8'd31;  //D
      
      //She said shut up.,...
      312: note<= 8'd31;  //D
	  313: note<= 8'd31;  //D
	  314: note<= 8'd25;  //Ab
      315: note<= 8'd25;  //Ab
      316: note<= 8'd23;  //F
      317: note<= 8'd21; //Eb
      318: note<= 8'd31;  //D
      319: note<= 8'd31;  //D
      
      //This woman is my ....
      320: note<= 8'd31;  //D
      321: note<= 8'd28; //Bb
      322: note<= 8'd31; //D
      323: note<= 8'd31; //D
      324: note<= 8'd21; //Eb
      325: note<= 8'd23; //F
      326: note<= 8'd31; //D
      327: note<= 8'd21; //Eb

//She siad ohh oh
      328: note<= 8'd31; //D
      329: note<= 8'd31; //D
      330: note<= 8'd25; //Ab
      331: note<= 8'd23; //F
      332: note<= 8'd28;  //Bb
      
      //Shut up and dance...
      333: note<= 8'd26; //Ab
      334: note<= 8'd26; //Ab
      335: note<= 8'd23; //F
      336: note<= 8'd21; //Eb
      337: note<= 8'd31;  //D
      338: note <= 8'd31;    //D
      */
    
	/*  0: note<= 8'd25;
	  1: note<= 8'd27;
	  2: note<= 8'd27;
	  3: note<= 8'd25;
	  4: note<= 8'd22;
	  5: note<= 8'd22;
	  6: note<= 8'd30;
	  7: note<= 8'd30;
	  8: note<= 8'd27;
	  9: note<= 8'd27;
	 10: note<= 8'd25;
	 11: note<= 8'd25;
	 12: note<= 8'd25;
	 13: note<= 8'd25;
	 14: note<= 8'd25;
	 15: note<= 8'd25;
	 16: note<= 8'd25;
	 17: note<= 8'd27;
	 18: note<= 8'd25;
	 19: note<= 8'd27;
	 20: note<= 8'd25;
	 21: note<= 8'd25;
	 22: note<= 8'd30;
	 23: note<= 8'd30;
	 24: note<= 8'd29;
	 25: note<= 8'd29;
	 26: note<= 8'd29;
	 27: note<= 8'd29;
	 28: note<= 8'd29;
	 29: note<= 8'd29;
	 30: note<= 8'd29;
	 31: note<= 8'd29;
	 32: note<= 8'd23;
	 33: note<= 8'd25;
	 34: note<= 8'd25;
	 35: note<= 8'd23;
	 36: note<= 8'd20;
	 37: note<= 8'd20;
	 38: note<= 8'd29;
	 39: note<= 8'd29;
	 40: note<= 8'd27;
	 41: note<= 8'd27;
	 42: note<= 8'd25;
	 43: note<= 8'd25;
	 44: note<= 8'd25;
	 45: note<= 8'd25;
	 46: note<= 8'd25;
	 47: note<= 8'd25;
	 48: note<= 8'd25;
	 49: note<= 8'd27;
	 50: note<= 8'd25;
	 51: note<= 8'd27;
	 52: note<= 8'd25;
	 53: note<= 8'd25;
	 54: note<= 8'd27;
	 55: note<= 8'd27;
	 56: note<= 8'd22;
	 57: note<= 8'd22;
	 58: note<= 8'd22;
	 59: note<= 8'd22;
	 60: note<= 8'd22;
	 61: note<= 8'd22;
	 62: note<= 8'd22;
	 63: note<= 8'd22;
	 64: note<= 8'd25;
	 65: note<= 8'd27;
	 66: note<= 8'd27;
	 67: note<= 8'd25;
	 68: note<= 8'd22;
	 69: note<= 8'd22;
	 70: note<= 8'd30;
	 71: note<= 8'd30;
	 72: note<= 8'd27;
	 73: note<= 8'd27;
	 74: note<= 8'd25;
	 75: note<= 8'd25;
	 76: note<= 8'd25;
	 77: note<= 8'd25;
	 78: note<= 8'd25;
	 79: note<= 8'd25;
	 80: note<= 8'd25;
	 81: note<= 8'd27;
	 82: note<= 8'd25;
	 83: note<= 8'd27;
	 84: note<= 8'd25;
	 85: note<= 8'd25;
	 86: note<= 8'd30;
	 87: note<= 8'd30;
	 88: note<= 8'd29;
	 89: note<= 8'd29;
	 90: note<= 8'd29;
	 91: note<= 8'd29;
	 92: note<= 8'd29;
	 93: note<= 8'd29;
	 94: note<= 8'd29;
	 95: note<= 8'd29;
	 96: note<= 8'd23;
	 97: note<= 8'd25;
	 98: note<= 8'd25;
	 99: note<= 8'd23;
	100: note<= 8'd20;
	101: note<= 8'd20;
	102: note<= 8'd29;
	103: note<= 8'd29;
	104: note<= 8'd27;
	105: note<= 8'd27;
	106: note<= 8'd25;
	107: note<= 8'd25;
	108: note<= 8'd25;
	109: note<= 8'd25;
	110: note<= 8'd25;
	111: note<= 8'd25;
	112: note<= 8'd25;
	113: note<= 8'd27;
	114: note<= 8'd25;
	115: note<= 8'd27;
	116: note<= 8'd25;
	117: note<= 8'd25;
	118: note<= 8'd32;
	119: note<= 8'd32;
	120: note<= 8'd30;
	121: note<= 8'd30;
	122: note<= 8'd30;
	123: note<= 8'd30;
	124: note<= 8'd30;
	125: note<= 8'd30;
	126: note<= 8'd30;
	127: note<= 8'd30;
	128: note<= 8'd27;
	129: note<= 8'd27;
	130: note<= 8'd27;
	131: note<= 8'd27;
	132: note<= 8'd30;
	133: note<= 8'd30;
	134: note<= 8'd30;
	135: note<= 8'd27;
	136: note<= 8'd25;
	137: note<= 8'd25;
	138: note<= 8'd22;
	139: note<= 8'd22;
	140: note<= 8'd25;
	141: note<= 8'd25;
	142: note<= 8'd25;
	143: note<= 8'd25;
	144: note<= 8'd23;
	145: note<= 8'd23;
	146: note<= 8'd27;
	147: note<= 8'd27;
	148: note<= 8'd25;
	149: note<= 8'd25;
	150: note<= 8'd23;
	151: note<= 8'd23;
	152: note<= 8'd22;
	153: note<= 8'd22;
	154: note<= 8'd22;
	155: note<= 8'd22;
	156: note<= 8'd22;
	157: note<= 8'd22;
	158: note<= 8'd22;
	159: note<= 8'd22;
	160: note<= 8'd20;
	161: note<= 8'd20;
	162: note<= 8'd22;
	163: note<= 8'd22;
	164: note<= 8'd25;
	165: note<= 8'd25;
	166: note<= 8'd27;
	167: note<= 8'd27;
	168: note<= 8'd29;
	169: note<= 8'd29;
	170: note<= 8'd29;
	171: note<= 8'd29;
	172: note<= 8'd29;
	173: note<= 8'd29;
	174: note<= 8'd29;
	175: note<= 8'd29;
	176: note<= 8'd30;
	177: note<= 8'd30;
	178: note<= 8'd30;
	179: note<= 8'd30;
	180: note<= 8'd29;
	181: note<= 8'd29;
	182: note<= 8'd27;
	183: note<= 8'd27;
	184: note<= 8'd25;
	185: note<= 8'd25;
	186: note<= 8'd23;
	187: note<= 8'd20;
	188: note<= 8'd20;
	189: note<= 8'd20;
	190: note<= 8'd20;
	191: note<= 8'd20;
	192: note<= 8'd25;
	193: note<= 8'd27;
	194: note<= 8'd27;
	195: note<= 8'd25;
	196: note<= 8'd22;
	197: note<= 8'd22;
	198: note<= 8'd30;
	199: note<= 8'd30;
	200: note<= 8'd27;
	201: note<= 8'd27;
	202: note<= 8'd25;
	203: note<= 8'd25;
	204: note<= 8'd25;
	205: note<= 8'd25;
	206: note<= 8'd25;
	207: note<= 8'd25;
	208: note<= 8'd25;
	209: note<= 8'd27;
	210: note<= 8'd25;
	211: note<= 8'd27;
	212: note<= 8'd25;
	213: note<= 8'd25;
	214: note<= 8'd30;
	215: note<= 8'd30;
	216: note<= 8'd29;
	217: note<= 8'd29;
	218: note<= 8'd29;
	219: note<= 8'd29;
	220: note<= 8'd29;
	221: note<= 8'd29;
	222: note<= 8'd29;
	223: note<= 8'd29;
	224: note<= 8'd23;
	225: note<= 8'd25;
	226: note<= 8'd25;
	227: note<= 8'd23;
	228: note<= 8'd20;
	229: note<= 8'd20;
	230: note<= 8'd29;
	231: note<= 8'd29;
	232: note<= 8'd27;
	233: note<= 8'd27;
	234: note<= 8'd25;
	235: note<= 8'd25;
	236: note<= 8'd25;
	237: note<= 8'd25;
	238: note<= 8'd25;
	239: note<= 8'd25;
	240: note<= 8'd25;
	241: note<= 8'd0;
	242: note<= 8'd00;*/

	default: note <= 8'd0;
endcase
endmodule